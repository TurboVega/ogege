/*
 * component_blender.v
 *
 * Copyright (C) 2024 by Curtis Whitley
 * License: APACHE
 */

`default_nettype none

module component_blender #(
) (
	input wire [3:0] i_bg_color,
	input wire [3:0] i_fg_color,
	input wire [2:0] i_fg_alpha,
	output wire [3:0] o_color
);

	wire [5:0] fg1 = {2'b0, i_fg_color};         // i_fg_color * 1, as 6 bits
	wire [5:0] fg2 = {1'b0, i_fg_color, 1'b0};   // i_fg_color * 2, as 6 bits
	wire [5:0] fg3 = fg1 + fg2;                  // i_fg_color * 3, as 6 bits

	wire [5:0] bg1 = {2'b0, i_bg_color};         // i_bg_color * 1, as 6 bits
	wire [5:0] bg2 = {1'b0, i_bg_color, 1'b0};   // i_bg_color * 2, as 6 bits
	wire [5:0] bg3 = bg1 + bg2;                  // i_bg_color * 3, as 6 bits

	wire [3:0] a;
	wire [3:0] b;
	wire [3:0] color;
	wire [5:0] sum;

	/*
		The "fg=33%, bg=67%" and "fg=67%, bg=33%" sub-case values below were generated by this code:

		#include <stdio.h>
		int main() {
			for (int a=0; a<16; a++) {
				for (int b=0; b<16; b++) {
					int c=(a+b*2)/3;
					printf("8'h%X%X: assign color = 4'h%X;\n",a,b,c);
				}
			}

			return 0;
		}
	*/

	case (i_fg_alpha)
		3'b000: assign color = i_bg_color;         	// fg=0%, bg=100%

		3'b001: begin								// fg=25%, bg=75%
					assign sum = (bg3 + fg1);
					assign color = sum[5:2];
				end

		3'b011: begin								// fg=50%, bg=50%
					assign sum = (bg1 + fg1);
					assign color = sum[4:1];
				end

		3'b101: begin								// fg=75%, bg=25%
					assign sum = (bg1 + fg3);
					assign color = sum[5:2];
				end

		3'b110: assign color = i_fg_color; 			// fg=100%, bg=0%

		3'b111: assign color = 4'b0000;              // reserved

		default: begin
			if (i_fg_alpha == 3'b010) begin
				// fg=33%, bg=67%
				assign a = i_fg_color;
				assign b = i_bg_color;
			end else begin // 3'b100
				// fg=67%, bg=33%
				assign a = i_bg_color;
				assign b = i_fg_color;
			end;

			case ({a, b})
				8'h00: assign color = 4'h0;
				8'h01: assign color = 4'h0;
				8'h02: assign color = 4'h1;
				8'h03: assign color = 4'h2;
				8'h04: assign color = 4'h2;
				8'h05: assign color = 4'h3;
				8'h06: assign color = 4'h4;
				8'h07: assign color = 4'h4;
				8'h08: assign color = 4'h5;
				8'h09: assign color = 4'h6;
				8'h0A: assign color = 4'h6;
				8'h0B: assign color = 4'h7;
				8'h0C: assign color = 4'h8;
				8'h0D: assign color = 4'h8;
				8'h0E: assign color = 4'h9;
				8'h0F: assign color = 4'hA;
				8'h10: assign color = 4'h0;
				8'h11: assign color = 4'h1;
				8'h12: assign color = 4'h1;
				8'h13: assign color = 4'h2;
				8'h14: assign color = 4'h3;
				8'h15: assign color = 4'h3;
				8'h16: assign color = 4'h4;
				8'h17: assign color = 4'h5;
				8'h18: assign color = 4'h5;
				8'h19: assign color = 4'h6;
				8'h1A: assign color = 4'h7;
				8'h1B: assign color = 4'h7;
				8'h1C: assign color = 4'h8;
				8'h1D: assign color = 4'h9;
				8'h1E: assign color = 4'h9;
				8'h1F: assign color = 4'hA;
				8'h20: assign color = 4'h0;
				8'h21: assign color = 4'h1;
				8'h22: assign color = 4'h2;
				8'h23: assign color = 4'h2;
				8'h24: assign color = 4'h3;
				8'h25: assign color = 4'h4;
				8'h26: assign color = 4'h4;
				8'h27: assign color = 4'h5;
				8'h28: assign color = 4'h6;
				8'h29: assign color = 4'h6;
				8'h2A: assign color = 4'h7;
				8'h2B: assign color = 4'h8;
				8'h2C: assign color = 4'h8;
				8'h2D: assign color = 4'h9;
				8'h2E: assign color = 4'hA;
				8'h2F: assign color = 4'hA;
				8'h30: assign color = 4'h1;
				8'h31: assign color = 4'h1;
				8'h32: assign color = 4'h2;
				8'h33: assign color = 4'h3;
				8'h34: assign color = 4'h3;
				8'h35: assign color = 4'h4;
				8'h36: assign color = 4'h5;
				8'h37: assign color = 4'h5;
				8'h38: assign color = 4'h6;
				8'h39: assign color = 4'h7;
				8'h3A: assign color = 4'h7;
				8'h3B: assign color = 4'h8;
				8'h3C: assign color = 4'h9;
				8'h3D: assign color = 4'h9;
				8'h3E: assign color = 4'hA;
				8'h3F: assign color = 4'hB;
				8'h40: assign color = 4'h1;
				8'h41: assign color = 4'h2;
				8'h42: assign color = 4'h2;
				8'h43: assign color = 4'h3;
				8'h44: assign color = 4'h4;
				8'h45: assign color = 4'h4;
				8'h46: assign color = 4'h5;
				8'h47: assign color = 4'h6;
				8'h48: assign color = 4'h6;
				8'h49: assign color = 4'h7;
				8'h4A: assign color = 4'h8;
				8'h4B: assign color = 4'h8;
				8'h4C: assign color = 4'h9;
				8'h4D: assign color = 4'hA;
				8'h4E: assign color = 4'hA;
				8'h4F: assign color = 4'hB;
				8'h50: assign color = 4'h1;
				8'h51: assign color = 4'h2;
				8'h52: assign color = 4'h3;
				8'h53: assign color = 4'h3;
				8'h54: assign color = 4'h4;
				8'h55: assign color = 4'h5;
				8'h56: assign color = 4'h5;
				8'h57: assign color = 4'h6;
				8'h58: assign color = 4'h7;
				8'h59: assign color = 4'h7;
				8'h5A: assign color = 4'h8;
				8'h5B: assign color = 4'h9;
				8'h5C: assign color = 4'h9;
				8'h5D: assign color = 4'hA;
				8'h5E: assign color = 4'hB;
				8'h5F: assign color = 4'hB;
				8'h60: assign color = 4'h2;
				8'h61: assign color = 4'h2;
				8'h62: assign color = 4'h3;
				8'h63: assign color = 4'h4;
				8'h64: assign color = 4'h4;
				8'h65: assign color = 4'h5;
				8'h66: assign color = 4'h6;
				8'h67: assign color = 4'h6;
				8'h68: assign color = 4'h7;
				8'h69: assign color = 4'h8;
				8'h6A: assign color = 4'h8;
				8'h6B: assign color = 4'h9;
				8'h6C: assign color = 4'hA;
				8'h6D: assign color = 4'hA;
				8'h6E: assign color = 4'hB;
				8'h6F: assign color = 4'hC;
				8'h70: assign color = 4'h2;
				8'h71: assign color = 4'h3;
				8'h72: assign color = 4'h3;
				8'h73: assign color = 4'h4;
				8'h74: assign color = 4'h5;
				8'h75: assign color = 4'h5;
				8'h76: assign color = 4'h6;
				8'h77: assign color = 4'h7;
				8'h78: assign color = 4'h7;
				8'h79: assign color = 4'h8;
				8'h7A: assign color = 4'h9;
				8'h7B: assign color = 4'h9;
				8'h7C: assign color = 4'hA;
				8'h7D: assign color = 4'hB;
				8'h7E: assign color = 4'hB;
				8'h7F: assign color = 4'hC;
				8'h80: assign color = 4'h2;
				8'h81: assign color = 4'h3;
				8'h82: assign color = 4'h4;
				8'h83: assign color = 4'h4;
				8'h84: assign color = 4'h5;
				8'h85: assign color = 4'h6;
				8'h86: assign color = 4'h6;
				8'h87: assign color = 4'h7;
				8'h88: assign color = 4'h8;
				8'h89: assign color = 4'h8;
				8'h8A: assign color = 4'h9;
				8'h8B: assign color = 4'hA;
				8'h8C: assign color = 4'hA;
				8'h8D: assign color = 4'hB;
				8'h8E: assign color = 4'hC;
				8'h8F: assign color = 4'hC;
				8'h90: assign color = 4'h3;
				8'h91: assign color = 4'h3;
				8'h92: assign color = 4'h4;
				8'h93: assign color = 4'h5;
				8'h94: assign color = 4'h5;
				8'h95: assign color = 4'h6;
				8'h96: assign color = 4'h7;
				8'h97: assign color = 4'h7;
				8'h98: assign color = 4'h8;
				8'h99: assign color = 4'h9;
				8'h9A: assign color = 4'h9;
				8'h9B: assign color = 4'hA;
				8'h9C: assign color = 4'hB;
				8'h9D: assign color = 4'hB;
				8'h9E: assign color = 4'hC;
				8'h9F: assign color = 4'hD;
				8'hA0: assign color = 4'h3;
				8'hA1: assign color = 4'h4;
				8'hA2: assign color = 4'h4;
				8'hA3: assign color = 4'h5;
				8'hA4: assign color = 4'h6;
				8'hA5: assign color = 4'h6;
				8'hA6: assign color = 4'h7;
				8'hA7: assign color = 4'h8;
				8'hA8: assign color = 4'h8;
				8'hA9: assign color = 4'h9;
				8'hAA: assign color = 4'hA;
				8'hAB: assign color = 4'hA;
				8'hAC: assign color = 4'hB;
				8'hAD: assign color = 4'hC;
				8'hAE: assign color = 4'hC;
				8'hAF: assign color = 4'hD;
				8'hB0: assign color = 4'h3;
				8'hB1: assign color = 4'h4;
				8'hB2: assign color = 4'h5;
				8'hB3: assign color = 4'h5;
				8'hB4: assign color = 4'h6;
				8'hB5: assign color = 4'h7;
				8'hB6: assign color = 4'h7;
				8'hB7: assign color = 4'h8;
				8'hB8: assign color = 4'h9;
				8'hB9: assign color = 4'h9;
				8'hBA: assign color = 4'hA;
				8'hBB: assign color = 4'hB;
				8'hBC: assign color = 4'hB;
				8'hBD: assign color = 4'hC;
				8'hBE: assign color = 4'hD;
				8'hBF: assign color = 4'hD;
				8'hC0: assign color = 4'h4;
				8'hC1: assign color = 4'h4;
				8'hC2: assign color = 4'h5;
				8'hC3: assign color = 4'h6;
				8'hC4: assign color = 4'h6;
				8'hC5: assign color = 4'h7;
				8'hC6: assign color = 4'h8;
				8'hC7: assign color = 4'h8;
				8'hC8: assign color = 4'h9;
				8'hC9: assign color = 4'hA;
				8'hCA: assign color = 4'hA;
				8'hCB: assign color = 4'hB;
				8'hCC: assign color = 4'hC;
				8'hCD: assign color = 4'hC;
				8'hCE: assign color = 4'hD;
				8'hCF: assign color = 4'hE;
				8'hD0: assign color = 4'h4;
				8'hD1: assign color = 4'h5;
				8'hD2: assign color = 4'h5;
				8'hD3: assign color = 4'h6;
				8'hD4: assign color = 4'h7;
				8'hD5: assign color = 4'h7;
				8'hD6: assign color = 4'h8;
				8'hD7: assign color = 4'h9;
				8'hD8: assign color = 4'h9;
				8'hD9: assign color = 4'hA;
				8'hDA: assign color = 4'hB;
				8'hDB: assign color = 4'hB;
				8'hDC: assign color = 4'hC;
				8'hDD: assign color = 4'hD;
				8'hDE: assign color = 4'hD;
				8'hDF: assign color = 4'hE;
				8'hE0: assign color = 4'h4;
				8'hE1: assign color = 4'h5;
				8'hE2: assign color = 4'h6;
				8'hE3: assign color = 4'h6;
				8'hE4: assign color = 4'h7;
				8'hE5: assign color = 4'h8;
				8'hE6: assign color = 4'h8;
				8'hE7: assign color = 4'h9;
				8'hE8: assign color = 4'hA;
				8'hE9: assign color = 4'hA;
				8'hEA: assign color = 4'hB;
				8'hEB: assign color = 4'hC;
				8'hEC: assign color = 4'hC;
				8'hED: assign color = 4'hD;
				8'hEE: assign color = 4'hE;
				8'hEF: assign color = 4'hE;
				8'hF0: assign color = 4'h5;
				8'hF1: assign color = 4'h5;
				8'hF2: assign color = 4'h6;
				8'hF3: assign color = 4'h7;
				8'hF4: assign color = 4'h7;
				8'hF5: assign color = 4'h8;
				8'hF6: assign color = 4'h9;
				8'hF7: assign color = 4'h9;
				8'hF8: assign color = 4'hA;
				8'hF9: assign color = 4'hB;
				8'hFA: assign color = 4'hB;
				8'hFB: assign color = 4'hC;
				8'hFC: assign color = 4'hD;
				8'hFD: assign color = 4'hD;
				8'hFE: assign color = 4'hE;
				8'hFF: assign color = 4'hF;
			endcase;
		end
	endcase;

	assign o_color = color;

endmodule
