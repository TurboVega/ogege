/*
 * component_blender.v
 *
 * Copyright (C) 2024 by Curtis Whitley
 * License: APACHE
 */

`default_nettype none

module component_blender #(
) (
	input wire [3:0] i_bg_color,
	input wire [3:0] i_fg_color,
	input wire [2:0] i_fg_alpha,
	output wire [3:0] o_color
);

	wire [5:0] fg1 = {2'b0, i_fg_color};         // i_fg_color * 1, as 6 bits
	wire [5:0] fg2 = {1'b0, i_fg_color, 1'b0};   // i_fg_color * 2, as 6 bits
	wire [5:0] fg3 = fg1 + fg2;                  // i_fg_color * 3, as 6 bits

	wire [5:0] bg1 = {2'b0, i_bg_color};         // i_bg_color * 1, as 6 bits
	wire [5:0] bg2 = {1'b0, i_bg_color, 1'b0};   // i_bg_color * 2, as 6 bits
	wire [5:0] bg3 = bg1 + bg2;                  // i_bg_color * 3, as 6 bits

	wire [3:0] a;
	wire [3:0] b;
	wire [3:0] color;

	/*
		The "fg=33%, bg=67%" and "fg=67%, bg=33%" sub-case values below were generated by this code:

		#include <stdio.h>
		int main() {
			for (int a=0; a<16; a++) {
				for (int b=0; b<16; b++) {
					int c=(a+b*2)/3;
					printf("8'h%X%X: color = 4'h%X;\n",a,b,c);
				}
			}

			return 0;
		}
	*/

	case (i_fg_alpha)
		3'b000: color = i_bg_color;           // fg=0%, bg=100%
		3'b001: color = (bg3 + fg1)[5:2];		// fg=25%, bg=75%
		3'b011: color = (bg1 + fg1)[4:1];		// fg=50%, bg=50%
		3'b101: color = (bg1 + fg3)[5:2];		// fg=75%, bg=25%
		3'b110: color = i_fg_color; 			// fg=100%, bg=0%
		3'b111: color = 4'b0000;              // reserved
		default: begin
			if (i_fg_alpha == 3'b010) begin
				// fg=33%, bg=67%
				a = i_fg_color;
				b = i_bg_color;
			end else begin // 3'b100
				// fg=67%, bg=33%
				a = i_bg_color;
				b = i_fg_color;
			end;

			case ({a, b})
				8'h00: color = 4'h0;
				8'h01: color = 4'h0;
				8'h02: color = 4'h1;
				8'h03: color = 4'h2;
				8'h04: color = 4'h2;
				8'h05: color = 4'h3;
				8'h06: color = 4'h4;
				8'h07: color = 4'h4;
				8'h08: color = 4'h5;
				8'h09: color = 4'h6;
				8'h0A: color = 4'h6;
				8'h0B: color = 4'h7;
				8'h0C: color = 4'h8;
				8'h0D: color = 4'h8;
				8'h0E: color = 4'h9;
				8'h0F: color = 4'hA;
				8'h10: color = 4'h0;
				8'h11: color = 4'h1;
				8'h12: color = 4'h1;
				8'h13: color = 4'h2;
				8'h14: color = 4'h3;
				8'h15: color = 4'h3;
				8'h16: color = 4'h4;
				8'h17: color = 4'h5;
				8'h18: color = 4'h5;
				8'h19: color = 4'h6;
				8'h1A: color = 4'h7;
				8'h1B: color = 4'h7;
				8'h1C: color = 4'h8;
				8'h1D: color = 4'h9;
				8'h1E: color = 4'h9;
				8'h1F: color = 4'hA;
				8'h20: color = 4'h0;
				8'h21: color = 4'h1;
				8'h22: color = 4'h2;
				8'h23: color = 4'h2;
				8'h24: color = 4'h3;
				8'h25: color = 4'h4;
				8'h26: color = 4'h4;
				8'h27: color = 4'h5;
				8'h28: color = 4'h6;
				8'h29: color = 4'h6;
				8'h2A: color = 4'h7;
				8'h2B: color = 4'h8;
				8'h2C: color = 4'h8;
				8'h2D: color = 4'h9;
				8'h2E: color = 4'hA;
				8'h2F: color = 4'hA;
				8'h30: color = 4'h1;
				8'h31: color = 4'h1;
				8'h32: color = 4'h2;
				8'h33: color = 4'h3;
				8'h34: color = 4'h3;
				8'h35: color = 4'h4;
				8'h36: color = 4'h5;
				8'h37: color = 4'h5;
				8'h38: color = 4'h6;
				8'h39: color = 4'h7;
				8'h3A: color = 4'h7;
				8'h3B: color = 4'h8;
				8'h3C: color = 4'h9;
				8'h3D: color = 4'h9;
				8'h3E: color = 4'hA;
				8'h3F: color = 4'hB;
				8'h40: color = 4'h1;
				8'h41: color = 4'h2;
				8'h42: color = 4'h2;
				8'h43: color = 4'h3;
				8'h44: color = 4'h4;
				8'h45: color = 4'h4;
				8'h46: color = 4'h5;
				8'h47: color = 4'h6;
				8'h48: color = 4'h6;
				8'h49: color = 4'h7;
				8'h4A: color = 4'h8;
				8'h4B: color = 4'h8;
				8'h4C: color = 4'h9;
				8'h4D: color = 4'hA;
				8'h4E: color = 4'hA;
				8'h4F: color = 4'hB;
				8'h50: color = 4'h1;
				8'h51: color = 4'h2;
				8'h52: color = 4'h3;
				8'h53: color = 4'h3;
				8'h54: color = 4'h4;
				8'h55: color = 4'h5;
				8'h56: color = 4'h5;
				8'h57: color = 4'h6;
				8'h58: color = 4'h7;
				8'h59: color = 4'h7;
				8'h5A: color = 4'h8;
				8'h5B: color = 4'h9;
				8'h5C: color = 4'h9;
				8'h5D: color = 4'hA;
				8'h5E: color = 4'hB;
				8'h5F: color = 4'hB;
				8'h60: color = 4'h2;
				8'h61: color = 4'h2;
				8'h62: color = 4'h3;
				8'h63: color = 4'h4;
				8'h64: color = 4'h4;
				8'h65: color = 4'h5;
				8'h66: color = 4'h6;
				8'h67: color = 4'h6;
				8'h68: color = 4'h7;
				8'h69: color = 4'h8;
				8'h6A: color = 4'h8;
				8'h6B: color = 4'h9;
				8'h6C: color = 4'hA;
				8'h6D: color = 4'hA;
				8'h6E: color = 4'hB;
				8'h6F: color = 4'hC;
				8'h70: color = 4'h2;
				8'h71: color = 4'h3;
				8'h72: color = 4'h3;
				8'h73: color = 4'h4;
				8'h74: color = 4'h5;
				8'h75: color = 4'h5;
				8'h76: color = 4'h6;
				8'h77: color = 4'h7;
				8'h78: color = 4'h7;
				8'h79: color = 4'h8;
				8'h7A: color = 4'h9;
				8'h7B: color = 4'h9;
				8'h7C: color = 4'hA;
				8'h7D: color = 4'hB;
				8'h7E: color = 4'hB;
				8'h7F: color = 4'hC;
				8'h80: color = 4'h2;
				8'h81: color = 4'h3;
				8'h82: color = 4'h4;
				8'h83: color = 4'h4;
				8'h84: color = 4'h5;
				8'h85: color = 4'h6;
				8'h86: color = 4'h6;
				8'h87: color = 4'h7;
				8'h88: color = 4'h8;
				8'h89: color = 4'h8;
				8'h8A: color = 4'h9;
				8'h8B: color = 4'hA;
				8'h8C: color = 4'hA;
				8'h8D: color = 4'hB;
				8'h8E: color = 4'hC;
				8'h8F: color = 4'hC;
				8'h90: color = 4'h3;
				8'h91: color = 4'h3;
				8'h92: color = 4'h4;
				8'h93: color = 4'h5;
				8'h94: color = 4'h5;
				8'h95: color = 4'h6;
				8'h96: color = 4'h7;
				8'h97: color = 4'h7;
				8'h98: color = 4'h8;
				8'h99: color = 4'h9;
				8'h9A: color = 4'h9;
				8'h9B: color = 4'hA;
				8'h9C: color = 4'hB;
				8'h9D: color = 4'hB;
				8'h9E: color = 4'hC;
				8'h9F: color = 4'hD;
				8'hA0: color = 4'h3;
				8'hA1: color = 4'h4;
				8'hA2: color = 4'h4;
				8'hA3: color = 4'h5;
				8'hA4: color = 4'h6;
				8'hA5: color = 4'h6;
				8'hA6: color = 4'h7;
				8'hA7: color = 4'h8;
				8'hA8: color = 4'h8;
				8'hA9: color = 4'h9;
				8'hAA: color = 4'hA;
				8'hAB: color = 4'hA;
				8'hAC: color = 4'hB;
				8'hAD: color = 4'hC;
				8'hAE: color = 4'hC;
				8'hAF: color = 4'hD;
				8'hB0: color = 4'h3;
				8'hB1: color = 4'h4;
				8'hB2: color = 4'h5;
				8'hB3: color = 4'h5;
				8'hB4: color = 4'h6;
				8'hB5: color = 4'h7;
				8'hB6: color = 4'h7;
				8'hB7: color = 4'h8;
				8'hB8: color = 4'h9;
				8'hB9: color = 4'h9;
				8'hBA: color = 4'hA;
				8'hBB: color = 4'hB;
				8'hBC: color = 4'hB;
				8'hBD: color = 4'hC;
				8'hBE: color = 4'hD;
				8'hBF: color = 4'hD;
				8'hC0: color = 4'h4;
				8'hC1: color = 4'h4;
				8'hC2: color = 4'h5;
				8'hC3: color = 4'h6;
				8'hC4: color = 4'h6;
				8'hC5: color = 4'h7;
				8'hC6: color = 4'h8;
				8'hC7: color = 4'h8;
				8'hC8: color = 4'h9;
				8'hC9: color = 4'hA;
				8'hCA: color = 4'hA;
				8'hCB: color = 4'hB;
				8'hCC: color = 4'hC;
				8'hCD: color = 4'hC;
				8'hCE: color = 4'hD;
				8'hCF: color = 4'hE;
				8'hD0: color = 4'h4;
				8'hD1: color = 4'h5;
				8'hD2: color = 4'h5;
				8'hD3: color = 4'h6;
				8'hD4: color = 4'h7;
				8'hD5: color = 4'h7;
				8'hD6: color = 4'h8;
				8'hD7: color = 4'h9;
				8'hD8: color = 4'h9;
				8'hD9: color = 4'hA;
				8'hDA: color = 4'hB;
				8'hDB: color = 4'hB;
				8'hDC: color = 4'hC;
				8'hDD: color = 4'hD;
				8'hDE: color = 4'hD;
				8'hDF: color = 4'hE;
				8'hE0: color = 4'h4;
				8'hE1: color = 4'h5;
				8'hE2: color = 4'h6;
				8'hE3: color = 4'h6;
				8'hE4: color = 4'h7;
				8'hE5: color = 4'h8;
				8'hE6: color = 4'h8;
				8'hE7: color = 4'h9;
				8'hE8: color = 4'hA;
				8'hE9: color = 4'hA;
				8'hEA: color = 4'hB;
				8'hEB: color = 4'hC;
				8'hEC: color = 4'hC;
				8'hED: color = 4'hD;
				8'hEE: color = 4'hE;
				8'hEF: color = 4'hE;
				8'hF0: color = 4'h5;
				8'hF1: color = 4'h5;
				8'hF2: color = 4'h6;
				8'hF3: color = 4'h7;
				8'hF4: color = 4'h7;
				8'hF5: color = 4'h8;
				8'hF6: color = 4'h9;
				8'hF7: color = 4'h9;
				8'hF8: color = 4'hA;
				8'hF9: color = 4'hB;
				8'hFA: color = 4'hB;
				8'hFB: color = 4'hC;
				8'hFC: color = 4'hD;
				8'hFD: color = 4'hD;
				8'hFE: color = 4'hE;
				8'hFF: color = 4'hF;
			endcase;
		end;
	endcase

	assign o_color = color;

endmodule
